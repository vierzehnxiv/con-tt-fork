/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_example (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  wire [31:0] lfsr_output;// = {16'b0, uio_out, uo_out};

  lfsr my_lfsr (
    .clk_i        (clk),
    .reset_i      (rst_n),
    .lfsr_state_o (lfsr_output) // only use lower 16 bits
  );

  // All output pins must be assigned. If not used, assign to 0.
  assign uio_oe  = 0;
  assign uio_out = lfsr_output[15:8];
  assign uo_out  = lfsr_output[7:0];
  //assign uo_out = 0;
  //assign uio_out = 0;

  // List all unused inputs to prevent warnings
  wire _unused = &{ui_in, uio_in, ena, 1'b0};

endmodule
